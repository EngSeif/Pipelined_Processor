--hello
--byeee
